module decrypt(clk,reset,data_in,data_out);
input clk;
input reset;
input [7:0] data_in;

output [7:0] data_out;

wire clk;
wire reset;
wire [7:0] data_in;

reg [7:0] data_out;

reg [7:0] mem [0:255];

always@(posedge clk)
    begin
      if(reset == 1)
          begin
         mem[0] <= 0;
         mem[1] <= 0;
         mem[2] <= 1;
         mem[3] <= 2;
         mem[4] <= 3;
         mem[5] <= 4;
         mem[6] <= 5;
         mem[7] <= 6;
         mem[8] <= 7;
         mem[9] <= 8;
         mem[10] <= 9;
         mem[11] <= 10;
         mem[12] <= 11;
         mem[13] <= 12;
         mem[14] <= 13;
         mem[15] <= 14;
         mem[16] <= 15;
         mem[17] <= 16;
         mem[18] <= 17;
         mem[19] <= 18;
         mem[20] <= 19;
         mem[21] <= 20;
         mem[22] <= 21;
         mem[23] <= 22;
         mem[24] <= 23;
         mem[25] <= 24;
         mem[26] <= 25;
         mem[27] <= 26;
         mem[28] <= 27;
         mem[29] <= 28;
         mem[30] <= 29;
         mem[31] <= 30;
         mem[32] <= 31;
         mem[33] <= 32;
         mem[34] <= 33;
         mem[35] <= 34;
         mem[36] <= 35;
         mem[37] <= 36;
         mem[38] <= 37;
         mem[39] <= 38;
         mem[40] <= 39;
         mem[41] <= 40;
         mem[42] <= 41;
         mem[43] <= 42;
         mem[44] <= 43;
         mem[45] <= 44;
         mem[46] <= 45;
         mem[47] <= 46;
         mem[48] <= 47;
         mem[49] <= 48;
         mem[50] <= 49;
         mem[51] <= 50;
         mem[52] <= 51;
         mem[53] <= 52;
         mem[54] <= 53;
         mem[55] <= 54;
         mem[56] <= 55;
         mem[57] <= 56;
         mem[58] <= 57;
         mem[59] <= 58;
         mem[60] <= 59;
         mem[61] <= 60;
         mem[62] <= 61;
         mem[63] <= 62;
         mem[64] <= 63;
         mem[65] <= 64;
         mem[66] <= 65;
         mem[67] <= 66;
         mem[68] <= 67;
         mem[69] <= 68;
         mem[70] <= 69;
         mem[71] <= 70;
         mem[72] <= 71;
         mem[73] <= 72;
         mem[74] <= 73;
         mem[75] <= 74;
         mem[76] <= 75;
         mem[77] <= 76;
         mem[78] <= 77;
         mem[79] <= 78;
         mem[80] <= 79;
         mem[81] <= 80;
         mem[82] <= 81;
         mem[83] <= 82;
         mem[84] <= 83;
         mem[85] <= 84;
         mem[86] <= 85;
         mem[87] <= 86;
         mem[88] <= 87;
         mem[89] <= 88;
         mem[90] <= 89;
         mem[91] <= 90;
         mem[92] <= 91;
         mem[93] <= 92;
         mem[94] <= 93;
         mem[95] <= 94;
         mem[96] <= 95;
         mem[97] <= 96;
         mem[98] <= 97;
         mem[99] <= 98;
         mem[100] <= 99;
         mem[101] <= 100;
         mem[102] <= 101;
         mem[103] <= 102;
         mem[104] <= 103;
         mem[105] <= 104;
         mem[106] <= 105;
         mem[107] <= 106;
         mem[108] <= 107;
         mem[109] <= 108;
         mem[110] <= 109;
         mem[111] <= 110;
         mem[112] <= 111;
         mem[113] <= 112;
         mem[114] <= 113;
         mem[115] <= 114;
         mem[116] <= 115;
         mem[117] <= 116;
         mem[118] <= 117;
         mem[119] <= 118;
         mem[120] <= 119;
         mem[121] <= 120;
         mem[122] <= 121;
         mem[123] <= 122;
         mem[124] <= 123;
         mem[125] <= 124;
         mem[126] <= 125;
         mem[127] <= 126;
         mem[128] <= 127;
         mem[129] <= 128;
         mem[130] <= 129;
         mem[131] <= 130;
         mem[132] <= 131;
         mem[133] <= 132;
         mem[134] <= 133;
         mem[135] <= 134;
         mem[136] <= 135;
         mem[137] <= 136;
         mem[138] <= 137;
         mem[139] <= 138;
         mem[140] <= 139;
         mem[141] <= 140;
         mem[142] <= 141;
         mem[143] <= 142;
         mem[144] <= 143;
         mem[145] <= 144;
         mem[146] <= 145;
         mem[147] <= 146;
         mem[148] <= 147;
         mem[149] <= 148;
         mem[150] <= 149;
         mem[151] <= 150;
         mem[152] <= 151;
         mem[153] <= 152;
         mem[154] <= 153;
         mem[155] <= 154;
         mem[156] <= 155;
         mem[157] <= 156;
         mem[158] <= 157;
         mem[159] <= 158;
         mem[160] <= 159;
         mem[161] <= 160;
         mem[162] <= 161;
         mem[163] <= 162;
         mem[164] <= 163;
         mem[165] <= 164;
         mem[166] <= 165;
         mem[167] <= 166;
         mem[168] <= 167;
         mem[169] <= 168;
         mem[170] <= 169;
         mem[171] <= 170;
         mem[172] <= 171;
         mem[173] <= 172;
         mem[174] <= 173;
         mem[175] <= 174;
         mem[176] <= 175;
         mem[177] <= 176;
         mem[178] <= 177;
         mem[179] <= 178;
         mem[180] <= 179;
         mem[181] <= 180;
         mem[182] <= 181;
         mem[183] <= 182;
         mem[184] <= 183;
         mem[185] <= 184;
         mem[186] <= 185;
         mem[187] <= 186;
         mem[188] <= 187;
         mem[189] <= 188;
         mem[190] <= 189;
         mem[191] <= 190;
         mem[192] <= 191;
         mem[193] <= 192;
         mem[194] <= 193;
         mem[195] <= 194;
         mem[196] <= 195;
         mem[197] <= 196;
         mem[198] <= 197;
         mem[199] <= 198;
         mem[200] <= 199;
         mem[201] <= 200;
         mem[202] <= 201;
         mem[203] <= 202;
         mem[204] <= 203;
         mem[205] <= 204;
         mem[206] <= 205;
         mem[207] <= 206;
         mem[208] <= 207;
         mem[209] <= 208;
         mem[210] <= 209;
         mem[211] <= 210;
         mem[212] <= 211;
         mem[213] <= 212;
         mem[214] <= 213;
         mem[215] <= 214;
         mem[216] <= 215;
         mem[217] <= 216;
         mem[218] <= 217;
         mem[219] <= 218;
         mem[220] <= 219;
         mem[221] <= 220;
         mem[222] <= 221;
         mem[223] <= 222;
         mem[224] <= 223;
         mem[225] <= 224;
         mem[226] <= 225;
         mem[227] <= 226;
         mem[228] <= 227;
         mem[229] <= 228;
         mem[230] <= 229;
         mem[231] <= 230;
         mem[232] <= 231;
         mem[233] <= 232;
         mem[234] <= 233;
         mem[235] <= 234;
         mem[236] <= 235;
         mem[237] <= 236;
         mem[238] <= 237;
         mem[239] <= 238;
         mem[240] <= 239;
         mem[241] <= 240;
         mem[242] <= 241;
         mem[243] <= 242;
         mem[244] <= 243;
         mem[245] <= 244;
         mem[246] <= 245;
         mem[247] <= 246;
         mem[248] <= 247;
         mem[249] <= 248;
         mem[250] <= 249;
         mem[251] <= 250;
         mem[252] <= 251;
         mem[253] <= 252;
         mem[254] <= 253;
         mem[255] <= 254;
         end
          else
            data_out <= mem[data_in];
end
endmodule
