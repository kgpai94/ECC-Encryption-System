module encrypt_y(clk,reset,data_in,data_out);
input clk;
input reset;
input [7:0] data_in;

output [7:0] data_out;

wire clk;
wire reset;
wire [7:0] data_in;

reg [7:0] data_out;

reg [7:0] mem [0:255];

always@(posedge clk)
begin
      if(reset == 1)
         begin
            mem[3] <= 8;
            mem[4] <= 3;
            mem[6] <= 8;
            mem[7] <= 5;
            mem[10] <= 6;
            mem[11] <= 8;
            mem[12] <= 7;
            mem[14] <= 11;
            mem[15] <= 6;
            mem[16] <= 1;
            mem[18] <= 6;
            mem[19] <= 7;
            mem[21] <= 2;
            mem[22] <= 2;
            mem[23] <= 2;
            mem[26] <= 8;
            mem[27] <= 3;
            mem[29] <= 8;
            mem[30] <= 5;
            mem[33] <= 6;
            mem[34] <= 8;
            mem[35] <= 7;
            mem[37] <= 11;
            mem[38] <= 6;
            mem[39] <= 1;
            mem[41] <= 6;
            mem[42] <= 7;
            mem[44] <= 2;
            mem[45] <= 2;
            mem[46] <= 2;
            mem[49] <= 8;
            mem[50] <= 3;
            mem[52] <= 8;
            mem[53] <= 5;
            mem[56] <= 6;
            mem[57] <= 8;
            mem[58] <= 7;
            mem[60] <= 11;
            mem[61] <= 6;
            mem[62] <= 1;
            mem[64] <= 6;
            mem[65] <= 7;
            mem[67] <= 2;
            mem[68] <= 2;
            mem[69] <= 2;
            mem[72] <= 8;
            mem[73] <= 3;
            mem[75] <= 8;
            mem[76] <= 5;
            mem[79] <= 6;
            mem[80] <= 8;
            mem[81] <= 7;
            mem[83] <= 11;
            mem[84] <= 6;
            mem[85] <= 1;
            mem[87] <= 6;
            mem[88] <= 7;
            mem[90] <= 2;
            mem[91] <= 2;
            mem[92] <= 2;
            mem[95] <= 8;
            mem[96] <= 3;
            mem[98] <= 8;
            mem[99] <= 5;
            mem[102] <= 6;
            mem[103] <= 8;
            mem[104] <= 7;
            mem[106] <= 11;
            mem[107] <= 6;
            mem[108] <= 1;
            mem[110] <= 6;
            mem[111] <= 7;
            mem[113] <= 2;
            mem[114] <= 2;
            mem[115] <= 2;
            mem[118] <= 8;
            mem[119] <= 3;
            mem[121] <= 8;
            mem[122] <= 5;
            mem[125] <= 6;
            mem[126] <= 8;
            mem[127] <= 7;
            mem[129] <= 11;
            mem[130] <= 6;
            mem[131] <= 1;
            mem[133] <= 6;
            mem[134] <= 7;
            mem[136] <= 2;
            mem[137] <= 2;
            mem[138] <= 2;
            mem[141] <= 8;
            mem[142] <= 3;
            mem[144] <= 8;
            mem[145] <= 5;
            mem[148] <= 6;
            mem[149] <= 8;
            mem[150] <= 7;
            mem[152] <= 11;
            mem[153] <= 6;
            mem[154] <= 1;
            mem[156] <= 6;
            mem[157] <= 7;
            mem[159] <= 2;
            mem[160] <= 2;
            mem[161] <= 2;
            mem[164] <= 8;
            mem[165] <= 3;
            mem[167] <= 8;
            mem[168] <= 5;
            mem[171] <= 6;
            mem[172] <= 8;
            mem[173] <= 7;
            mem[175] <= 11;
            mem[176] <= 6;
            mem[177] <= 1;
            mem[179] <= 6;
            mem[180] <= 7;
            mem[182] <= 2;
            mem[183] <= 2;
            mem[184] <= 2;
            mem[187] <= 8;
            mem[188] <= 3;
            mem[190] <= 8;
            mem[191] <= 5;
            mem[194] <= 6;
            mem[195] <= 8;
            mem[196] <= 7;
            mem[198] <= 11;
            mem[199] <= 6;
            mem[200] <= 1;
            mem[202] <= 6;
            mem[203] <= 7;
            mem[205] <= 2;
            mem[206] <= 2;
            mem[207] <= 2;
            mem[210] <= 8;
            mem[211] <= 3;
            mem[213] <= 8;
            mem[214] <= 5;
            mem[217] <= 6;
            mem[218] <= 8;
            mem[219] <= 7;
            mem[221] <= 11;
            mem[222] <= 6;
            mem[223] <= 1;
            mem[225] <= 6;
            mem[226] <= 7;
            mem[228] <= 2;
            mem[229] <= 2;
            mem[230] <= 2;
            mem[233] <= 8;
            mem[234] <= 3;
            mem[236] <= 8;
            mem[237] <= 5;
            mem[240] <= 6;
            mem[241] <= 8;
            mem[242] <= 7;
            mem[244] <= 11;
            mem[245] <= 6;
            mem[246] <= 1;
            mem[248] <= 6;
            mem[249] <= 7;
            mem[251] <= 2;
            mem[252] <= 2;
            mem[253] <= 2;
          end

          else
              data_out <= mem[data_in];

  end

endmodule  
